magic
tech sky130A
magscale 1 2
timestamp 1716990733
<< locali >>
rect 15572 42186 15616 42196
rect 15572 42152 15577 42186
rect 15611 42152 15616 42186
rect 15572 42114 15616 42152
rect 15572 42080 15577 42114
rect 15611 42080 15616 42114
rect 15572 42042 15616 42080
rect 15572 42008 15577 42042
rect 15611 42008 15616 42042
rect 15572 41970 15616 42008
rect 15572 41936 15577 41970
rect 15611 41936 15616 41970
rect 14756 41888 15144 41932
rect 15572 41898 15616 41936
rect 15572 41864 15577 41898
rect 15611 41864 15616 41898
rect 15572 41826 15616 41864
rect 15572 41792 15577 41826
rect 15611 41792 15616 41826
rect 15572 41754 15616 41792
rect 15572 41720 15577 41754
rect 15611 41720 15616 41754
rect 15572 41682 15616 41720
rect 15572 41648 15577 41682
rect 15611 41648 15616 41682
rect 15572 41610 15616 41648
rect 15572 41576 15577 41610
rect 15611 41576 15616 41610
rect 15572 41538 15616 41576
rect 15572 41504 15577 41538
rect 15611 41504 15616 41538
rect 15572 41466 15616 41504
rect 15572 41432 15577 41466
rect 15611 41432 15616 41466
rect 18218 42191 18264 42192
rect 18218 42157 18224 42191
rect 18258 42157 18264 42191
rect 21220 42174 21266 42196
rect 18218 42119 18264 42157
rect 18218 42085 18224 42119
rect 18258 42085 18264 42119
rect 18218 42047 18264 42085
rect 18218 42013 18224 42047
rect 18258 42013 18264 42047
rect 18218 41975 18264 42013
rect 18218 41941 18224 41975
rect 18258 41941 18264 41975
rect 18218 41903 18264 41941
rect 18218 41869 18224 41903
rect 18258 41869 18264 41903
rect 18670 42158 18714 42168
rect 18670 42124 18675 42158
rect 18709 42124 18714 42158
rect 18670 42086 18714 42124
rect 18670 42052 18675 42086
rect 18709 42052 18714 42086
rect 18670 42014 18714 42052
rect 18670 41980 18675 42014
rect 18709 41980 18714 42014
rect 18670 41942 18714 41980
rect 18670 41908 18675 41942
rect 18709 41908 18714 41942
rect 18670 41898 18714 41908
rect 19956 42158 20004 42168
rect 19956 42124 19963 42158
rect 19997 42124 20004 42158
rect 19956 42086 20004 42124
rect 19956 42052 19963 42086
rect 19997 42052 20004 42086
rect 19956 42014 20004 42052
rect 19956 41980 19963 42014
rect 19997 41980 20004 42014
rect 19956 41942 20004 41980
rect 19956 41908 19963 41942
rect 19997 41908 20004 41942
rect 19956 41898 20004 41908
rect 21220 42140 21226 42174
rect 21260 42140 21266 42174
rect 21220 42102 21266 42140
rect 21220 42068 21226 42102
rect 21260 42068 21266 42102
rect 21220 42030 21266 42068
rect 21220 41996 21226 42030
rect 21260 41996 21266 42030
rect 21220 41958 21266 41996
rect 21220 41924 21226 41958
rect 21260 41924 21266 41958
rect 21220 41902 21266 41924
rect 21744 41890 22132 41932
rect 18218 41831 18264 41869
rect 18218 41797 18224 41831
rect 18258 41797 18264 41831
rect 18218 41759 18264 41797
rect 18218 41725 18224 41759
rect 18258 41725 18264 41759
rect 18218 41687 18264 41725
rect 18218 41653 18224 41687
rect 18258 41653 18264 41687
rect 18218 41615 18264 41653
rect 18218 41581 18224 41615
rect 18258 41581 18264 41615
rect 18218 41543 18264 41581
rect 18218 41509 18224 41543
rect 18258 41509 18264 41543
rect 18218 41471 18264 41509
rect 18218 41437 18224 41471
rect 18258 41437 18264 41471
rect 18218 41436 18264 41437
rect 15572 41422 15616 41432
rect 20330 41370 20376 41380
rect 20330 41336 20336 41370
rect 20370 41336 20376 41370
rect 20330 41298 20376 41336
rect 20330 41264 20336 41298
rect 20370 41264 20376 41298
rect 20330 41226 20376 41264
rect 20330 41192 20336 41226
rect 20370 41192 20376 41226
rect 20330 41154 20376 41192
rect 20330 41120 20336 41154
rect 20370 41120 20376 41154
rect 20330 41082 20376 41120
rect 20330 41048 20336 41082
rect 20370 41048 20376 41082
rect 20330 41010 20376 41048
rect 20330 40976 20336 41010
rect 20370 40976 20376 41010
rect 20330 40938 20376 40976
rect 20330 40904 20336 40938
rect 20370 40904 20376 40938
rect 15574 40893 15618 40904
rect 15574 40859 15579 40893
rect 15613 40859 15618 40893
rect 15574 40821 15618 40859
rect 15574 40787 15579 40821
rect 15613 40787 15618 40821
rect 15574 40749 15618 40787
rect 15574 40715 15579 40749
rect 15613 40715 15618 40749
rect 15574 40677 15618 40715
rect 15574 40643 15579 40677
rect 15613 40643 15618 40677
rect 15574 40605 15618 40643
rect 15574 40571 15579 40605
rect 15613 40571 15618 40605
rect 15574 40533 15618 40571
rect 15574 40499 15579 40533
rect 15613 40499 15618 40533
rect 15574 40461 15618 40499
rect 15574 40427 15579 40461
rect 15613 40427 15618 40461
rect 15574 40389 15618 40427
rect 15574 40355 15579 40389
rect 15613 40355 15618 40389
rect 15574 40317 15618 40355
rect 15574 40283 15579 40317
rect 15613 40283 15618 40317
rect 15574 40245 15618 40283
rect 15574 40211 15579 40245
rect 15613 40211 15618 40245
rect 15574 40173 15618 40211
rect 15574 40139 15579 40173
rect 15613 40139 15618 40173
rect 15574 40128 15618 40139
rect 16462 40893 16504 40904
rect 16462 40859 16466 40893
rect 16500 40859 16504 40893
rect 16462 40821 16504 40859
rect 16462 40787 16466 40821
rect 16500 40787 16504 40821
rect 16462 40749 16504 40787
rect 16462 40715 16466 40749
rect 16500 40715 16504 40749
rect 16462 40677 16504 40715
rect 16462 40643 16466 40677
rect 16500 40643 16504 40677
rect 16462 40605 16504 40643
rect 20330 40866 20376 40904
rect 20330 40832 20336 40866
rect 20370 40832 20376 40866
rect 20330 40794 20376 40832
rect 20330 40760 20336 40794
rect 20370 40760 20376 40794
rect 20330 40722 20376 40760
rect 20330 40688 20336 40722
rect 20370 40688 20376 40722
rect 20330 40650 20376 40688
rect 20330 40616 20336 40650
rect 20370 40616 20376 40650
rect 20330 40606 20376 40616
rect 21216 41370 21262 41380
rect 21216 41336 21222 41370
rect 21256 41336 21262 41370
rect 21216 41298 21262 41336
rect 21216 41264 21222 41298
rect 21256 41264 21262 41298
rect 21216 41226 21262 41264
rect 21216 41192 21222 41226
rect 21256 41192 21262 41226
rect 21216 41154 21262 41192
rect 21216 41120 21222 41154
rect 21256 41120 21262 41154
rect 21216 41082 21262 41120
rect 21216 41048 21222 41082
rect 21256 41048 21262 41082
rect 21216 41010 21262 41048
rect 21216 40976 21222 41010
rect 21256 40976 21262 41010
rect 21216 40938 21262 40976
rect 21216 40904 21222 40938
rect 21256 40904 21262 40938
rect 21216 40866 21262 40904
rect 21216 40832 21222 40866
rect 21256 40832 21262 40866
rect 21216 40794 21262 40832
rect 21216 40760 21222 40794
rect 21256 40760 21262 40794
rect 21216 40722 21262 40760
rect 21216 40688 21222 40722
rect 21256 40688 21262 40722
rect 21216 40650 21262 40688
rect 21216 40616 21222 40650
rect 21256 40616 21262 40650
rect 21216 40606 21262 40616
rect 16462 40571 16466 40605
rect 16500 40571 16504 40605
rect 16462 40533 16504 40571
rect 16462 40499 16466 40533
rect 16500 40499 16504 40533
rect 16462 40461 16504 40499
rect 16462 40427 16466 40461
rect 16500 40427 16504 40461
rect 16462 40389 16504 40427
rect 16462 40355 16466 40389
rect 16500 40355 16504 40389
rect 16462 40317 16504 40355
rect 16462 40283 16466 40317
rect 16500 40283 16504 40317
rect 16462 40245 16504 40283
rect 16462 40211 16466 40245
rect 16500 40211 16504 40245
rect 16462 40173 16504 40211
rect 16462 40139 16466 40173
rect 16500 40139 16504 40173
rect 16462 40128 16504 40139
rect 20332 40076 20378 40086
rect 18668 40065 18712 40066
rect 18668 40031 18673 40065
rect 18707 40031 18712 40065
rect 18668 39993 18712 40031
rect 18668 39959 18673 39993
rect 18707 39959 18712 39993
rect 18668 39921 18712 39959
rect 18668 39887 18673 39921
rect 18707 39887 18712 39921
rect 18668 39849 18712 39887
rect 18668 39815 18673 39849
rect 18707 39815 18712 39849
rect 18668 39777 18712 39815
rect 18668 39743 18673 39777
rect 18707 39743 18712 39777
rect 18668 39705 18712 39743
rect 18668 39671 18673 39705
rect 18707 39671 18712 39705
rect 18668 39633 18712 39671
rect 15572 39586 15616 39608
rect 15572 39552 15577 39586
rect 15611 39552 15616 39586
rect 15572 39514 15616 39552
rect 15572 39480 15577 39514
rect 15611 39480 15616 39514
rect 15572 39442 15616 39480
rect 15572 39408 15577 39442
rect 15611 39408 15616 39442
rect 15572 39370 15616 39408
rect 15572 39336 15577 39370
rect 15611 39336 15616 39370
rect 15572 39314 15616 39336
rect 16458 39586 16502 39608
rect 16458 39552 16463 39586
rect 16497 39552 16502 39586
rect 18668 39599 18673 39633
rect 18707 39599 18712 39633
rect 16458 39514 16502 39552
rect 16458 39480 16463 39514
rect 16497 39480 16502 39514
rect 16458 39442 16502 39480
rect 16458 39408 16463 39442
rect 16497 39408 16502 39442
rect 16458 39370 16502 39408
rect 16458 39336 16463 39370
rect 16497 39336 16502 39370
rect 16458 39314 16502 39336
rect 16858 39572 16910 39582
rect 16858 39538 16867 39572
rect 16901 39538 16910 39572
rect 16858 39500 16910 39538
rect 16858 39466 16867 39500
rect 16901 39466 16910 39500
rect 16858 39428 16910 39466
rect 16858 39394 16867 39428
rect 16901 39394 16910 39428
rect 16858 39356 16910 39394
rect 16858 39322 16867 39356
rect 16901 39322 16910 39356
rect 16858 39312 16910 39322
rect 18148 39572 18196 39582
rect 18148 39538 18155 39572
rect 18189 39538 18196 39572
rect 18148 39500 18196 39538
rect 18148 39466 18155 39500
rect 18189 39466 18196 39500
rect 18148 39428 18196 39466
rect 18148 39394 18155 39428
rect 18189 39394 18196 39428
rect 18148 39356 18196 39394
rect 18148 39322 18155 39356
rect 18189 39322 18196 39356
rect 18148 39312 18196 39322
rect 18668 39561 18712 39599
rect 18668 39527 18673 39561
rect 18707 39527 18712 39561
rect 18668 39489 18712 39527
rect 18668 39455 18673 39489
rect 18707 39455 18712 39489
rect 18668 39417 18712 39455
rect 18668 39383 18673 39417
rect 18707 39383 18712 39417
rect 18668 39345 18712 39383
rect 18668 39311 18673 39345
rect 18707 39311 18712 39345
rect 20332 40042 20338 40076
rect 20372 40042 20378 40076
rect 20332 40004 20378 40042
rect 20332 39970 20338 40004
rect 20372 39970 20378 40004
rect 20332 39932 20378 39970
rect 20332 39898 20338 39932
rect 20372 39898 20378 39932
rect 20332 39860 20378 39898
rect 20332 39826 20338 39860
rect 20372 39826 20378 39860
rect 20332 39788 20378 39826
rect 20332 39754 20338 39788
rect 20372 39754 20378 39788
rect 20332 39716 20378 39754
rect 20332 39682 20338 39716
rect 20372 39682 20378 39716
rect 20332 39644 20378 39682
rect 20332 39610 20338 39644
rect 20372 39610 20378 39644
rect 20332 39572 20378 39610
rect 20332 39538 20338 39572
rect 20372 39538 20378 39572
rect 20332 39500 20378 39538
rect 20332 39466 20338 39500
rect 20372 39466 20378 39500
rect 20332 39428 20378 39466
rect 20332 39394 20338 39428
rect 20372 39394 20378 39428
rect 20332 39356 20378 39394
rect 20332 39322 20338 39356
rect 20372 39322 20378 39356
rect 20332 39312 20378 39322
rect 21220 40076 21262 40086
rect 21220 40042 21224 40076
rect 21258 40042 21262 40076
rect 21220 40004 21262 40042
rect 21220 39970 21224 40004
rect 21258 39970 21262 40004
rect 21220 39932 21262 39970
rect 21220 39898 21224 39932
rect 21258 39898 21262 39932
rect 21220 39860 21262 39898
rect 21220 39826 21224 39860
rect 21258 39826 21262 39860
rect 21220 39788 21262 39826
rect 21220 39754 21224 39788
rect 21258 39754 21262 39788
rect 21220 39716 21262 39754
rect 21220 39682 21224 39716
rect 21258 39682 21262 39716
rect 21220 39644 21262 39682
rect 21220 39610 21224 39644
rect 21258 39610 21262 39644
rect 21220 39572 21262 39610
rect 21220 39538 21224 39572
rect 21258 39538 21262 39572
rect 21220 39500 21262 39538
rect 21220 39466 21224 39500
rect 21258 39466 21262 39500
rect 21220 39428 21262 39466
rect 21220 39394 21224 39428
rect 21258 39394 21262 39428
rect 21220 39356 21262 39394
rect 21220 39322 21224 39356
rect 21258 39322 21262 39356
rect 21220 39312 21262 39322
rect 18668 39310 18712 39311
<< viali >>
rect 15577 42152 15611 42186
rect 15577 42080 15611 42114
rect 15577 42008 15611 42042
rect 15577 41936 15611 41970
rect 15577 41864 15611 41898
rect 15577 41792 15611 41826
rect 15577 41720 15611 41754
rect 15577 41648 15611 41682
rect 15577 41576 15611 41610
rect 15577 41504 15611 41538
rect 15577 41432 15611 41466
rect 18224 42157 18258 42191
rect 18224 42085 18258 42119
rect 18224 42013 18258 42047
rect 18224 41941 18258 41975
rect 18224 41869 18258 41903
rect 18675 42124 18709 42158
rect 18675 42052 18709 42086
rect 18675 41980 18709 42014
rect 18675 41908 18709 41942
rect 19963 42124 19997 42158
rect 19963 42052 19997 42086
rect 19963 41980 19997 42014
rect 19963 41908 19997 41942
rect 21226 42140 21260 42174
rect 21226 42068 21260 42102
rect 21226 41996 21260 42030
rect 21226 41924 21260 41958
rect 18224 41797 18258 41831
rect 18224 41725 18258 41759
rect 18224 41653 18258 41687
rect 18224 41581 18258 41615
rect 18224 41509 18258 41543
rect 18224 41437 18258 41471
rect 20336 41336 20370 41370
rect 20336 41264 20370 41298
rect 20336 41192 20370 41226
rect 20336 41120 20370 41154
rect 20336 41048 20370 41082
rect 20336 40976 20370 41010
rect 20336 40904 20370 40938
rect 15579 40859 15613 40893
rect 15579 40787 15613 40821
rect 15579 40715 15613 40749
rect 15579 40643 15613 40677
rect 15579 40571 15613 40605
rect 15579 40499 15613 40533
rect 15579 40427 15613 40461
rect 15579 40355 15613 40389
rect 15579 40283 15613 40317
rect 15579 40211 15613 40245
rect 15579 40139 15613 40173
rect 16466 40859 16500 40893
rect 16466 40787 16500 40821
rect 16466 40715 16500 40749
rect 16466 40643 16500 40677
rect 20336 40832 20370 40866
rect 20336 40760 20370 40794
rect 20336 40688 20370 40722
rect 20336 40616 20370 40650
rect 21222 41336 21256 41370
rect 21222 41264 21256 41298
rect 21222 41192 21256 41226
rect 21222 41120 21256 41154
rect 21222 41048 21256 41082
rect 21222 40976 21256 41010
rect 21222 40904 21256 40938
rect 21222 40832 21256 40866
rect 21222 40760 21256 40794
rect 21222 40688 21256 40722
rect 21222 40616 21256 40650
rect 16466 40571 16500 40605
rect 16466 40499 16500 40533
rect 16466 40427 16500 40461
rect 16466 40355 16500 40389
rect 16466 40283 16500 40317
rect 16466 40211 16500 40245
rect 16466 40139 16500 40173
rect 18673 40031 18707 40065
rect 18673 39959 18707 39993
rect 18673 39887 18707 39921
rect 18673 39815 18707 39849
rect 18673 39743 18707 39777
rect 18673 39671 18707 39705
rect 15577 39552 15611 39586
rect 15577 39480 15611 39514
rect 15577 39408 15611 39442
rect 15577 39336 15611 39370
rect 16463 39552 16497 39586
rect 18673 39599 18707 39633
rect 16463 39480 16497 39514
rect 16463 39408 16497 39442
rect 16463 39336 16497 39370
rect 16867 39538 16901 39572
rect 16867 39466 16901 39500
rect 16867 39394 16901 39428
rect 16867 39322 16901 39356
rect 18155 39538 18189 39572
rect 18155 39466 18189 39500
rect 18155 39394 18189 39428
rect 18155 39322 18189 39356
rect 18673 39527 18707 39561
rect 18673 39455 18707 39489
rect 18673 39383 18707 39417
rect 18673 39311 18707 39345
rect 20338 40042 20372 40076
rect 20338 39970 20372 40004
rect 20338 39898 20372 39932
rect 20338 39826 20372 39860
rect 20338 39754 20372 39788
rect 20338 39682 20372 39716
rect 20338 39610 20372 39644
rect 20338 39538 20372 39572
rect 20338 39466 20372 39500
rect 20338 39394 20372 39428
rect 20338 39322 20372 39356
rect 21224 40042 21258 40076
rect 21224 39970 21258 40004
rect 21224 39898 21258 39932
rect 21224 39826 21258 39860
rect 21224 39754 21258 39788
rect 21224 39682 21258 39716
rect 21224 39610 21258 39644
rect 21224 39538 21258 39572
rect 21224 39466 21258 39500
rect 21224 39394 21258 39428
rect 21224 39322 21258 39356
<< metal1 >>
rect 14373 42830 23529 42841
rect 14373 42778 23470 42830
rect 23522 42778 23529 42830
rect 14373 42767 23529 42778
rect 14373 42345 14447 42767
rect 14608 42632 21316 42652
rect 14608 42580 14672 42632
rect 14724 42580 21316 42632
rect 14608 42560 21316 42580
rect 14373 42271 14747 42345
rect 15572 42304 15620 42560
rect 19862 42396 20474 42434
rect 14673 41950 14747 42271
rect 15560 42186 15630 42304
rect 15560 42152 15577 42186
rect 15611 42152 15630 42186
rect 15560 42114 15630 42152
rect 15560 42080 15577 42114
rect 15611 42080 15630 42114
rect 15560 42042 15630 42080
rect 18210 42191 18280 42308
rect 18210 42157 18224 42191
rect 18258 42157 18280 42191
rect 18210 42119 18280 42157
rect 18210 42085 18224 42119
rect 18258 42085 18280 42119
rect 18210 42052 18280 42085
rect 18658 42158 18728 42280
rect 18658 42124 18675 42158
rect 18709 42124 18728 42158
rect 18658 42086 18728 42124
rect 18658 42052 18675 42086
rect 18709 42052 18728 42086
rect 19862 42072 19906 42396
rect 19944 42158 20020 42282
rect 19944 42124 19963 42158
rect 19997 42124 20020 42158
rect 19944 42086 20020 42124
rect 19944 42052 19963 42086
rect 19997 42052 20020 42086
rect 20430 42072 20474 42396
rect 21226 42308 21274 42560
rect 21208 42174 21282 42308
rect 21208 42140 21226 42174
rect 21260 42140 21282 42174
rect 21208 42102 21282 42140
rect 21208 42068 21226 42102
rect 21260 42068 21282 42102
rect 21208 42062 21282 42068
rect 15560 42008 15577 42042
rect 15611 42008 15630 42042
rect 15560 41970 15630 42008
rect 18130 42047 18802 42052
rect 18130 42013 18224 42047
rect 18258 42014 18802 42047
rect 18258 42013 18675 42014
rect 18130 41990 18675 42013
rect 14648 41874 15258 41950
rect 15560 41936 15577 41970
rect 15611 41936 15630 41970
rect 15560 41898 15630 41936
rect 15560 41864 15577 41898
rect 15611 41864 15630 41898
rect 15560 41834 15630 41864
rect 18210 41975 18280 41990
rect 18210 41941 18224 41975
rect 18258 41941 18280 41975
rect 18210 41903 18280 41941
rect 18210 41869 18224 41903
rect 18258 41869 18280 41903
rect 14772 41740 14832 41828
rect 15560 41826 15722 41834
rect 15560 41792 15577 41826
rect 15611 41792 15722 41826
rect 16366 41794 17070 41846
rect 18210 41831 18280 41869
rect 18210 41797 18224 41831
rect 18258 41797 18280 41831
rect 15560 41788 15722 41792
rect 15560 41754 15630 41788
rect 15560 41720 15577 41754
rect 15611 41720 15630 41754
rect 15560 41682 15630 41720
rect 15560 41648 15577 41682
rect 15611 41648 15630 41682
rect 15560 41610 15630 41648
rect 15560 41576 15577 41610
rect 15611 41576 15630 41610
rect 15560 41538 15630 41576
rect 18210 41759 18280 41797
rect 18658 41980 18675 41990
rect 18709 41990 18802 42014
rect 19944 42014 20020 42052
rect 21120 42030 21282 42062
rect 21120 42020 21226 42030
rect 18709 41980 18728 41990
rect 18658 41942 18728 41980
rect 19944 41980 19963 42014
rect 19997 41980 20020 42014
rect 18658 41908 18675 41942
rect 18709 41908 18728 41942
rect 18658 41788 18728 41908
rect 18210 41725 18224 41759
rect 18258 41725 18280 41759
rect 18210 41687 18280 41725
rect 18210 41653 18224 41687
rect 18258 41653 18280 41687
rect 18210 41615 18280 41653
rect 18210 41581 18224 41615
rect 18258 41581 18280 41615
rect 15560 41504 15577 41538
rect 15611 41504 15630 41538
rect 15560 41466 15630 41504
rect 15560 41432 15577 41466
rect 15611 41432 15630 41466
rect 15560 40893 15630 41432
rect 15560 40859 15579 40893
rect 15613 40859 15630 40893
rect 15996 40882 16056 41458
rect 17064 41438 17132 41558
rect 18210 41543 18280 41581
rect 18210 41509 18224 41543
rect 18258 41509 18280 41543
rect 18210 41471 18280 41509
rect 17988 41198 18056 41466
rect 18210 41437 18224 41471
rect 18258 41437 18280 41471
rect 18210 41328 18280 41437
rect 18876 41198 18948 41950
rect 19944 41942 20020 41980
rect 19944 41908 19963 41942
rect 19997 41908 20020 41942
rect 21208 41996 21226 42020
rect 21260 41996 21282 42030
rect 21208 41958 21282 41996
rect 19944 41786 20020 41908
rect 17988 41124 18948 41198
rect 17988 41122 18056 41124
rect 15560 40821 15630 40859
rect 15560 40787 15579 40821
rect 15613 40787 15630 40821
rect 15560 40749 15630 40787
rect 16322 40768 16388 40900
rect 16450 40893 16514 41022
rect 16450 40859 16466 40893
rect 16500 40859 16514 40893
rect 16450 40821 16514 40859
rect 16450 40787 16466 40821
rect 16500 40787 16514 40821
rect 15560 40715 15579 40749
rect 15613 40715 15630 40749
rect 15560 40677 15630 40715
rect 15560 40643 15579 40677
rect 15613 40643 15630 40677
rect 15560 40605 15630 40643
rect 15560 40571 15579 40605
rect 15613 40571 15630 40605
rect 15560 40534 15630 40571
rect 16450 40749 16514 40787
rect 19954 40784 20008 41786
rect 16450 40715 16466 40749
rect 16500 40715 16514 40749
rect 16450 40677 16514 40715
rect 16450 40643 16466 40677
rect 16500 40643 16514 40677
rect 16450 40605 16514 40643
rect 16450 40571 16466 40605
rect 16500 40571 16514 40605
rect 15560 40533 15718 40534
rect 15560 40499 15579 40533
rect 15613 40499 15718 40533
rect 15560 40490 15718 40499
rect 16450 40533 16514 40571
rect 16450 40499 16466 40533
rect 16500 40499 16514 40533
rect 15560 40461 15630 40490
rect 15560 40427 15579 40461
rect 15613 40427 15630 40461
rect 15560 40389 15630 40427
rect 15560 40355 15579 40389
rect 15613 40355 15630 40389
rect 15560 40317 15630 40355
rect 15560 40283 15579 40317
rect 15613 40283 15630 40317
rect 15560 40245 15630 40283
rect 15560 40211 15579 40245
rect 15613 40211 15630 40245
rect 15560 40173 15630 40211
rect 15560 40139 15579 40173
rect 15613 40139 15630 40173
rect 16450 40461 16514 40499
rect 16450 40427 16466 40461
rect 16500 40427 16514 40461
rect 16450 40389 16514 40427
rect 16450 40355 16466 40389
rect 16500 40355 16514 40389
rect 16450 40317 16514 40355
rect 16450 40283 16466 40317
rect 16500 40283 16514 40317
rect 16450 40245 16514 40283
rect 16450 40211 16466 40245
rect 16500 40211 16514 40245
rect 16450 40173 16514 40211
rect 15560 40022 15630 40139
rect 15996 39870 16056 40152
rect 15110 39818 16056 39870
rect 14754 38966 14794 39776
rect 15560 39586 15630 39714
rect 15560 39552 15577 39586
rect 15611 39552 15630 39586
rect 15996 39576 16056 39818
rect 16450 40139 16466 40173
rect 16500 40139 16514 40173
rect 16450 39586 16514 40139
rect 16852 40716 20008 40784
rect 20320 41370 20392 41496
rect 20320 41336 20336 41370
rect 20370 41336 20392 41370
rect 20738 41362 20798 41938
rect 21208 41924 21226 41958
rect 21260 41924 21282 41958
rect 22132 42267 23508 42278
rect 22132 42215 23431 42267
rect 23483 42215 23508 42267
rect 22132 42206 23508 42215
rect 22132 41942 22204 42206
rect 21208 41370 21282 41924
rect 21632 41870 22242 41942
rect 22058 41734 22118 41822
rect 20320 41298 20392 41336
rect 20320 41264 20336 41298
rect 20370 41264 20392 41298
rect 20320 41226 20392 41264
rect 20320 41192 20336 41226
rect 20370 41192 20392 41226
rect 20320 41154 20392 41192
rect 20320 41120 20336 41154
rect 20370 41120 20392 41154
rect 20320 41082 20392 41120
rect 20320 41048 20336 41082
rect 20370 41048 20392 41082
rect 20320 41010 20392 41048
rect 20320 40976 20336 41010
rect 20370 40976 20392 41010
rect 21208 41336 21222 41370
rect 21256 41336 21282 41370
rect 21208 41298 21282 41336
rect 21208 41264 21222 41298
rect 21256 41264 21282 41298
rect 21208 41226 21282 41264
rect 21208 41192 21222 41226
rect 21256 41192 21282 41226
rect 21208 41154 21282 41192
rect 21208 41120 21222 41154
rect 21256 41120 21282 41154
rect 21208 41082 21282 41120
rect 21208 41048 21222 41082
rect 21256 41048 21282 41082
rect 21208 41010 21282 41048
rect 21208 41008 21222 41010
rect 20320 40938 20392 40976
rect 21116 40976 21222 41008
rect 21256 40976 21282 41010
rect 21116 40968 21282 40976
rect 20320 40904 20336 40938
rect 20370 40904 20392 40938
rect 20320 40866 20392 40904
rect 20320 40832 20336 40866
rect 20370 40832 20392 40866
rect 20320 40794 20392 40832
rect 20320 40760 20336 40794
rect 20370 40760 20392 40794
rect 20320 40722 20392 40760
rect 21208 40938 21282 40968
rect 21208 40904 21222 40938
rect 21256 40904 21282 40938
rect 21208 40866 21282 40904
rect 21208 40832 21222 40866
rect 21256 40832 21282 40866
rect 21208 40794 21282 40832
rect 21208 40760 21222 40794
rect 21256 40760 21282 40794
rect 16852 39694 16916 40716
rect 20320 40688 20336 40722
rect 20370 40688 20392 40722
rect 20320 40650 20392 40688
rect 20320 40616 20336 40650
rect 20370 40616 20392 40650
rect 20452 40616 20518 40748
rect 21208 40722 21282 40760
rect 21208 40688 21222 40722
rect 21256 40688 21282 40722
rect 21208 40650 21282 40688
rect 17976 40308 18936 40382
rect 15560 39514 15630 39552
rect 15560 39480 15577 39514
rect 15611 39482 15630 39514
rect 16450 39552 16463 39586
rect 16497 39552 16514 39586
rect 16450 39514 16514 39552
rect 15611 39480 15712 39482
rect 15560 39442 15712 39480
rect 16450 39480 16463 39514
rect 16497 39480 16514 39514
rect 15560 39408 15577 39442
rect 15611 39440 15712 39442
rect 15611 39408 15630 39440
rect 15560 39370 15630 39408
rect 15560 39336 15577 39370
rect 15611 39336 15630 39370
rect 15560 39210 15630 39336
rect 16362 39148 16410 39462
rect 16450 39442 16514 39480
rect 16450 39408 16463 39442
rect 16497 39408 16514 39442
rect 16450 39370 16514 39408
rect 16450 39336 16463 39370
rect 16497 39336 16514 39370
rect 16450 39200 16514 39336
rect 16842 39572 16920 39694
rect 16842 39538 16867 39572
rect 16901 39538 16920 39572
rect 17976 39556 18048 40308
rect 18656 40065 18720 40184
rect 18656 40031 18673 40065
rect 18707 40031 18720 40065
rect 18868 40038 18936 40308
rect 20320 40076 20392 40616
rect 18656 39993 18720 40031
rect 18656 39959 18673 39993
rect 18707 39959 18720 39993
rect 19808 39966 19876 40064
rect 20320 40042 20338 40076
rect 20372 40042 20392 40076
rect 20808 40352 20868 40638
rect 21208 40616 21222 40650
rect 21256 40616 21282 40650
rect 21208 40492 21282 40616
rect 20808 40300 21786 40352
rect 20808 40062 20868 40300
rect 21210 40076 21278 40198
rect 20320 40004 20392 40042
rect 20320 39970 20338 40004
rect 20372 39970 20392 40004
rect 18656 39921 18720 39959
rect 18656 39887 18673 39921
rect 18707 39887 18720 39921
rect 18656 39849 18720 39887
rect 18656 39815 18673 39849
rect 18707 39815 18720 39849
rect 18656 39777 18720 39815
rect 18656 39743 18673 39777
rect 18707 39743 18720 39777
rect 18656 39705 18720 39743
rect 18140 39572 18214 39694
rect 16842 39500 16920 39538
rect 16842 39466 16867 39500
rect 16901 39466 16920 39500
rect 18140 39538 18155 39572
rect 18189 39538 18214 39572
rect 18140 39500 18214 39538
rect 18140 39484 18155 39500
rect 16842 39428 16920 39466
rect 18058 39466 18155 39484
rect 18189 39484 18214 39500
rect 18656 39671 18673 39705
rect 18707 39671 18720 39705
rect 18656 39633 18720 39671
rect 18656 39599 18673 39633
rect 18707 39599 18720 39633
rect 18656 39561 18720 39599
rect 18656 39527 18673 39561
rect 18707 39527 18720 39561
rect 18656 39489 18720 39527
rect 18656 39484 18673 39489
rect 18189 39466 18673 39484
rect 16842 39394 16867 39428
rect 16901 39394 16920 39428
rect 16842 39356 16920 39394
rect 16842 39322 16867 39356
rect 16901 39322 16920 39356
rect 16842 39202 16920 39322
rect 16952 39148 17000 39462
rect 18058 39455 18673 39466
rect 18707 39484 18720 39489
rect 20320 39932 20392 39970
rect 20320 39898 20338 39932
rect 20372 39898 20392 39932
rect 20320 39860 20392 39898
rect 20320 39826 20338 39860
rect 20372 39826 20392 39860
rect 20320 39788 20392 39826
rect 20320 39754 20338 39788
rect 20372 39754 20392 39788
rect 20320 39716 20392 39754
rect 21210 40042 21224 40076
rect 21258 40042 21278 40076
rect 21210 40004 21278 40042
rect 21210 39970 21224 40004
rect 21258 39970 21278 40004
rect 21210 39932 21278 39970
rect 21210 39898 21224 39932
rect 21258 39898 21278 39932
rect 21210 39860 21278 39898
rect 21210 39826 21224 39860
rect 21258 39826 21278 39860
rect 21210 39788 21278 39826
rect 21210 39754 21224 39788
rect 21258 39754 21278 39788
rect 21210 39718 21278 39754
rect 20320 39682 20338 39716
rect 20372 39682 20392 39716
rect 20320 39644 20392 39682
rect 21118 39716 21278 39718
rect 21118 39682 21224 39716
rect 21258 39682 21278 39716
rect 21118 39678 21278 39682
rect 20320 39610 20338 39644
rect 20372 39610 20392 39644
rect 20320 39572 20392 39610
rect 20320 39538 20338 39572
rect 20372 39538 20392 39572
rect 20320 39500 20392 39538
rect 18707 39455 18806 39484
rect 18058 39428 18806 39455
rect 20320 39466 20338 39500
rect 20372 39466 20392 39500
rect 18058 39422 18155 39428
rect 18140 39394 18155 39422
rect 18189 39422 18806 39428
rect 18189 39394 18214 39422
rect 18140 39356 18214 39394
rect 18140 39322 18155 39356
rect 18189 39322 18214 39356
rect 18140 39200 18214 39322
rect 16362 39096 17000 39148
rect 16714 39082 16798 39096
rect 16714 39030 16729 39082
rect 16781 39030 16798 39082
rect 16714 39018 16798 39030
rect 18360 38966 18452 39422
rect 18656 39417 18720 39422
rect 18656 39383 18673 39417
rect 18707 39383 18720 39417
rect 18656 39345 18720 39383
rect 18656 39311 18673 39345
rect 18707 39311 18720 39345
rect 18656 39202 18720 39311
rect 19876 39144 19920 39438
rect 20320 39428 20392 39466
rect 21210 39644 21278 39678
rect 21210 39610 21224 39644
rect 21258 39610 21278 39644
rect 21210 39572 21278 39610
rect 21210 39538 21224 39572
rect 21258 39538 21278 39572
rect 21210 39500 21278 39538
rect 21210 39466 21224 39500
rect 21258 39466 21278 39500
rect 20320 39394 20338 39428
rect 20372 39394 20392 39428
rect 20320 39356 20392 39394
rect 20320 39322 20338 39356
rect 20372 39322 20392 39356
rect 20320 39200 20392 39322
rect 20428 39144 20472 39438
rect 21210 39428 21278 39466
rect 21210 39394 21224 39428
rect 21258 39394 21278 39428
rect 21210 39356 21278 39394
rect 21210 39322 21224 39356
rect 21258 39322 21278 39356
rect 21210 39198 21278 39322
rect 19876 39092 20472 39144
rect 22098 38966 22138 39778
rect 14632 38937 22262 38966
rect 14632 38885 15011 38937
rect 15063 38885 22262 38937
rect 14632 38860 22262 38885
<< via1 >>
rect 23470 42778 23522 42830
rect 14672 42580 14724 42632
rect 23431 42215 23483 42267
rect 16729 39030 16781 39082
rect 15011 38885 15063 38937
<< metal2 >>
rect 23448 42833 23540 42846
rect 23448 42777 23463 42833
rect 23519 42830 23540 42833
rect 23522 42778 23540 42830
rect 23519 42777 23540 42778
rect 23448 42762 23540 42777
rect 8145 42639 14774 42696
rect 8145 42583 8282 42639
rect 8338 42632 14774 42639
rect 8338 42583 14672 42632
rect 8145 42580 14672 42583
rect 14724 42580 14774 42632
rect 8145 42522 14774 42580
rect 23406 42270 23508 42284
rect 23406 42214 23429 42270
rect 23485 42214 23508 42270
rect 23406 42196 23508 42214
rect 16704 39085 16818 39108
rect 16704 39029 16727 39085
rect 16783 39029 16818 39085
rect 16704 39010 16818 39029
rect 14958 38941 15116 38988
rect 14958 38885 15008 38941
rect 15064 38885 15116 38941
rect 14958 38834 15116 38885
<< via2 >>
rect 23463 42830 23519 42833
rect 23463 42778 23470 42830
rect 23470 42778 23519 42830
rect 23463 42777 23519 42778
rect 8282 42583 8338 42639
rect 23429 42267 23485 42270
rect 23429 42215 23431 42267
rect 23431 42215 23483 42267
rect 23483 42215 23485 42267
rect 23429 42214 23485 42215
rect 16727 39082 16783 39085
rect 16727 39030 16729 39082
rect 16729 39030 16781 39082
rect 16781 39030 16783 39082
rect 16727 39029 16783 39030
rect 15008 38937 15064 38941
rect 15008 38885 15011 38937
rect 15011 38885 15063 38937
rect 15063 38885 15064 38937
<< metal3 >>
rect 23440 42837 23552 42862
rect 23440 42773 23457 42837
rect 23521 42773 23552 42837
rect 23440 42756 23552 42773
rect 8140 42641 8458 42716
rect 8140 42577 8238 42641
rect 8302 42639 8318 42641
rect 8302 42577 8318 42583
rect 8382 42577 8458 42641
rect 8140 42496 8458 42577
rect 23422 42274 23492 42278
rect 23422 42210 23425 42274
rect 23489 42210 23492 42274
rect 23422 42206 23492 42210
rect 16698 39089 16824 39112
rect 16698 39025 16723 39089
rect 16787 39025 16824 39089
rect 16698 39006 16824 39025
rect 14940 38942 15136 39004
rect 14940 38878 15005 38942
rect 15069 38878 15136 38942
rect 14940 38814 15136 38878
<< rmetal3 >>
rect 23400 42278 23514 42290
rect 23400 42206 23422 42278
rect 23492 42206 23514 42278
rect 23400 42190 23514 42206
<< via3 >>
rect 23457 42833 23521 42837
rect 23457 42777 23463 42833
rect 23463 42777 23519 42833
rect 23519 42777 23521 42833
rect 23457 42773 23521 42777
rect 8238 42639 8302 42641
rect 8318 42639 8382 42641
rect 8238 42583 8282 42639
rect 8282 42583 8302 42639
rect 8318 42583 8338 42639
rect 8338 42583 8382 42639
rect 8238 42577 8302 42583
rect 8318 42577 8382 42583
rect 23425 42270 23489 42274
rect 23425 42214 23429 42270
rect 23429 42214 23485 42270
rect 23485 42214 23489 42270
rect 23425 42210 23489 42214
rect 16723 39085 16787 39089
rect 16723 39029 16727 39085
rect 16727 39029 16783 39085
rect 16783 39029 16787 39085
rect 16723 39025 16787 39029
rect 15005 38941 15069 38942
rect 15005 38885 15008 38941
rect 15008 38885 15064 38941
rect 15064 38885 15069 38941
rect 15005 38878 15069 38885
<< metal4 >>
rect 798 45092 858 45152
rect 1534 45092 1594 45152
rect 2270 45092 2330 45152
rect 3006 45092 3066 45152
rect 3742 45092 3802 45152
rect 4478 45092 4538 45152
rect 5214 45092 5274 45152
rect 5950 45092 6010 45152
rect 6686 45092 6746 45152
rect 7422 45092 7482 45152
rect 8158 45092 8218 45152
rect 8894 45092 8954 45152
rect 9630 45092 9690 45152
rect 10366 45092 10426 45152
rect 11102 45092 11162 45152
rect 11838 45092 11898 45152
rect 12574 45092 12634 45152
rect 13310 45092 13370 45152
rect 14046 45092 14106 45152
rect 14782 45092 14842 45152
rect 15518 45092 15578 45152
rect 16254 45092 16314 45152
rect 16990 45092 17050 45152
rect 17726 45092 17786 45152
rect 798 44974 17786 45092
rect 798 44952 858 44974
rect 1534 44952 1594 44974
rect 2270 44952 2330 44974
rect 3006 44952 3066 44974
rect 3742 44952 3802 44974
rect 4478 44952 4538 44974
rect 5214 44952 5274 44974
rect 5950 44952 6010 44974
rect 6686 44952 6746 44974
rect 7422 44952 7482 44974
rect 8158 44952 8218 44974
rect 8894 44952 8954 44974
rect 9630 44952 9690 44974
rect 10366 44952 10426 44974
rect 11102 44952 11162 44974
rect 11838 44952 11898 44974
rect 200 42770 500 44152
rect 200 42641 8494 42770
rect 200 42577 8238 42641
rect 8302 42577 8318 42641
rect 8382 42577 8494 42641
rect 200 42470 8494 42577
rect 200 1000 500 42470
rect 9800 39050 10100 44152
rect 12533 39050 12651 44974
rect 13310 44952 13370 44974
rect 14046 44952 14106 44974
rect 14782 44952 14842 44974
rect 15518 44952 15578 44974
rect 16254 44952 16314 44974
rect 16990 44950 17050 44974
rect 17726 44950 17786 44974
rect 18462 44952 18522 45152
rect 19198 44952 19258 45152
rect 19934 44952 19994 45152
rect 20670 44952 20730 45152
rect 21406 44952 21466 45152
rect 22142 44952 22202 45152
rect 22878 44952 22938 45152
rect 23614 44952 23674 45152
rect 24350 44952 24410 45152
rect 25086 44952 25146 45152
rect 25822 44952 25882 45152
rect 26558 44952 26618 45152
rect 27294 44952 27354 45152
rect 28030 44952 28090 45152
rect 28766 44952 28826 45152
rect 29502 44948 29562 45152
rect 30238 44952 30298 45152
rect 30974 44952 31034 45152
rect 31710 44952 31770 45152
rect 23348 42837 31462 42896
rect 23348 42773 23457 42837
rect 23521 42773 31462 42837
rect 23348 42716 31462 42773
rect 23380 42274 27046 42332
rect 23380 42210 23425 42274
rect 23489 42210 27046 42274
rect 23380 42152 27046 42210
rect 16678 39089 16846 39128
rect 9800 38942 15198 39050
rect 9800 38878 15005 38942
rect 15069 38878 15198 38942
rect 9800 38750 15198 38878
rect 16678 39025 16723 39089
rect 16787 39025 16846 39089
rect 9800 1000 10100 38750
rect 16678 38300 16846 39025
rect 16678 38120 22630 38300
rect 370 0 550 200
rect 4786 0 4966 200
rect 9202 0 9382 200
rect 13618 0 13798 200
rect 18034 0 18214 200
rect 22450 0 22630 38120
rect 26866 0 27046 42152
rect 31282 0 31462 42716
use sky130_fd_pr__nfet_01v8_HXU4AK  sky130_fd_pr__nfet_01v8_HXU4AK_0
timestamp 1716990733
transform 1 0 19336 0 1 42033
box -686 -257 686 257
use sky130_fd_pr__nfet_01v8_HXU4AK  sky130_fd_pr__nfet_01v8_HXU4AK_1
timestamp 1716990733
transform 1 0 17528 0 1 39447
box -686 -257 686 257
use sky130_fd_pr__nfet_01v8_MXF53G  sky130_fd_pr__nfet_01v8_MXF53G_0
timestamp 1716990733
transform 1 0 19332 0 1 39688
box -686 -500 686 500
use sky130_fd_pr__nfet_01v8_MXF53G  sky130_fd_pr__nfet_01v8_MXF53G_1
timestamp 1716990733
transform 1 0 17598 0 1 41814
box -686 -500 686 500
use sky130_fd_pr__pfet_01v8_GE7BQD  sky130_fd_pr__pfet_01v8_GE7BQD_0
timestamp 1716990733
transform 1 0 14950 0 1 40745
box -326 -1219 326 1219
use sky130_fd_pr__pfet_01v8_GE7BQD  sky130_fd_pr__pfet_01v8_GE7BQD_1
timestamp 1716990733
transform 1 0 21938 0 1 40745
box -326 -1219 326 1219
use sky130_fd_pr__pfet_01v8_KDYT8F  sky130_fd_pr__pfet_01v8_KDYT8F_0
timestamp 1716990733
transform 1 0 20800 0 1 42049
box -496 -279 496 279
use sky130_fd_pr__pfet_01v8_KDYT8F  sky130_fd_pr__pfet_01v8_KDYT8F_1
timestamp 1716990733
transform 1 0 16036 0 1 39461
box -496 -279 496 279
use sky130_fd_pr__pfet_01v8_NXK9QA  sky130_fd_pr__pfet_01v8_NXK9QA_0
timestamp 1716990733
transform -1 0 16039 0 -1 40516
box -496 -519 496 519
use sky130_fd_pr__pfet_01v8_NXK9QA  sky130_fd_pr__pfet_01v8_NXK9QA_1
timestamp 1716990733
transform -1 0 20798 0 -1 39699
box -496 -519 496 519
use sky130_fd_pr__pfet_01v8_NXK9QA  sky130_fd_pr__pfet_01v8_NXK9QA_2
timestamp 1716990733
transform -1 0 16038 0 -1 41809
box -496 -519 496 519
use sky130_fd_pr__pfet_01v8_NXK9QA  sky130_fd_pr__pfet_01v8_NXK9QA_3
timestamp 1716990733
transform -1 0 20796 0 -1 40993
box -496 -519 496 519
<< labels >>
flabel metal4 s 30974 44952 31034 45152 0 FreeSans 600 90 0 0 clk
flabel metal4 s 31710 44952 31770 45152 0 FreeSans 600 90 0 0 ena
flabel metal4 s 30238 44952 30298 45152 0 FreeSans 600 90 0 0 rst_n
flabel metal4 s 31282 0 31462 200 0 FreeSans 1200 0 0 0 ua[0]
flabel metal4 s 26866 0 27046 200 0 FreeSans 1200 0 0 0 ua[1]
flabel metal4 s 22450 0 22630 200 0 FreeSans 1200 0 0 0 ua[2]
flabel metal4 s 18034 0 18214 200 0 FreeSans 1200 0 0 0 ua[3]
flabel metal4 s 13618 0 13798 200 0 FreeSans 1200 0 0 0 ua[4]
flabel metal4 s 9202 0 9382 200 0 FreeSans 1200 0 0 0 ua[5]
flabel metal4 s 4786 0 4966 200 0 FreeSans 1200 0 0 0 ua[6]
flabel metal4 s 370 0 550 200 0 FreeSans 1200 0 0 0 ua[7]
flabel metal4 s 29502 44952 29562 45152 0 FreeSans 600 90 0 0 ui_in[0]
flabel metal4 s 28766 44952 28826 45152 0 FreeSans 600 90 0 0 ui_in[1]
flabel metal4 s 28030 44952 28090 45152 0 FreeSans 600 90 0 0 ui_in[2]
flabel metal4 s 27294 44952 27354 45152 0 FreeSans 600 90 0 0 ui_in[3]
flabel metal4 s 26558 44952 26618 45152 0 FreeSans 600 90 0 0 ui_in[4]
flabel metal4 s 25822 44952 25882 45152 0 FreeSans 600 90 0 0 ui_in[5]
flabel metal4 s 25086 44952 25146 45152 0 FreeSans 600 90 0 0 ui_in[6]
flabel metal4 s 24350 44952 24410 45152 0 FreeSans 600 90 0 0 ui_in[7]
flabel metal4 s 23614 44952 23674 45152 0 FreeSans 600 90 0 0 uio_in[0]
flabel metal4 s 22878 44952 22938 45152 0 FreeSans 600 90 0 0 uio_in[1]
flabel metal4 s 22142 44952 22202 45152 0 FreeSans 600 90 0 0 uio_in[2]
flabel metal4 s 21406 44952 21466 45152 0 FreeSans 600 90 0 0 uio_in[3]
flabel metal4 s 20670 44952 20730 45152 0 FreeSans 600 90 0 0 uio_in[4]
flabel metal4 s 19934 44952 19994 45152 0 FreeSans 600 90 0 0 uio_in[5]
flabel metal4 s 19198 44952 19258 45152 0 FreeSans 600 90 0 0 uio_in[6]
flabel metal4 s 18462 44952 18522 45152 0 FreeSans 600 90 0 0 uio_in[7]
flabel metal4 s 5950 44952 6010 45152 0 FreeSans 600 90 0 0 uio_oe[0]
flabel metal4 s 5214 44952 5274 45152 0 FreeSans 600 90 0 0 uio_oe[1]
flabel metal4 s 4478 44952 4538 45152 0 FreeSans 600 90 0 0 uio_oe[2]
flabel metal4 s 3742 44952 3802 45152 0 FreeSans 600 90 0 0 uio_oe[3]
flabel metal4 s 3006 44952 3066 45152 0 FreeSans 600 90 0 0 uio_oe[4]
flabel metal4 s 2270 44952 2330 45152 0 FreeSans 600 90 0 0 uio_oe[5]
flabel metal4 s 1534 44952 1594 45152 0 FreeSans 600 90 0 0 uio_oe[6]
flabel metal4 s 798 44952 858 45152 0 FreeSans 600 90 0 0 uio_oe[7]
flabel metal4 s 11838 44952 11898 45152 0 FreeSans 600 90 0 0 uio_out[0]
flabel metal4 s 11102 44952 11162 45152 0 FreeSans 600 90 0 0 uio_out[1]
flabel metal4 s 10366 44952 10426 45152 0 FreeSans 600 90 0 0 uio_out[2]
flabel metal4 s 9630 44952 9690 45152 0 FreeSans 600 90 0 0 uio_out[3]
flabel metal4 s 8894 44952 8954 45152 0 FreeSans 600 90 0 0 uio_out[4]
flabel metal4 s 8158 44952 8218 45152 0 FreeSans 600 90 0 0 uio_out[5]
flabel metal4 s 7422 44952 7482 45152 0 FreeSans 600 90 0 0 uio_out[6]
flabel metal4 s 6686 44952 6746 45152 0 FreeSans 600 90 0 0 uio_out[7]
flabel metal4 s 17726 44952 17786 45152 0 FreeSans 600 90 0 0 uo_out[0]
flabel metal4 s 16990 44952 17050 45152 0 FreeSans 600 90 0 0 uo_out[1]
flabel metal4 s 16254 44952 16314 45152 0 FreeSans 600 90 0 0 uo_out[2]
flabel metal4 s 15518 44952 15578 45152 0 FreeSans 600 90 0 0 uo_out[3]
flabel metal4 s 14782 44952 14842 45152 0 FreeSans 600 90 0 0 uo_out[4]
flabel metal4 s 14046 44952 14106 45152 0 FreeSans 600 90 0 0 uo_out[5]
flabel metal4 s 13310 44952 13370 45152 0 FreeSans 600 90 0 0 uo_out[6]
flabel metal4 s 12574 44952 12634 45152 0 FreeSans 600 90 0 0 uo_out[7]
flabel metal4 s 200 1000 500 44152 1 FreeSans 2 0 0 0 VPWR
flabel metal4 s 9800 1000 10100 44152 1 FreeSans 2 0 0 0 VGND
<< properties >>
string FIXED_BBOX 0 0 32200 45152
<< end >>
