magic
tech sky130A
magscale 1 2
timestamp 1716990733
<< nwell >>
rect -326 -1219 326 1219
<< pmos >>
rect -130 -1000 130 1000
<< pdiff >>
rect -188 969 -130 1000
rect -188 935 -176 969
rect -142 935 -130 969
rect -188 901 -130 935
rect -188 867 -176 901
rect -142 867 -130 901
rect -188 833 -130 867
rect -188 799 -176 833
rect -142 799 -130 833
rect -188 765 -130 799
rect -188 731 -176 765
rect -142 731 -130 765
rect -188 697 -130 731
rect -188 663 -176 697
rect -142 663 -130 697
rect -188 629 -130 663
rect -188 595 -176 629
rect -142 595 -130 629
rect -188 561 -130 595
rect -188 527 -176 561
rect -142 527 -130 561
rect -188 493 -130 527
rect -188 459 -176 493
rect -142 459 -130 493
rect -188 425 -130 459
rect -188 391 -176 425
rect -142 391 -130 425
rect -188 357 -130 391
rect -188 323 -176 357
rect -142 323 -130 357
rect -188 289 -130 323
rect -188 255 -176 289
rect -142 255 -130 289
rect -188 221 -130 255
rect -188 187 -176 221
rect -142 187 -130 221
rect -188 153 -130 187
rect -188 119 -176 153
rect -142 119 -130 153
rect -188 85 -130 119
rect -188 51 -176 85
rect -142 51 -130 85
rect -188 17 -130 51
rect -188 -17 -176 17
rect -142 -17 -130 17
rect -188 -51 -130 -17
rect -188 -85 -176 -51
rect -142 -85 -130 -51
rect -188 -119 -130 -85
rect -188 -153 -176 -119
rect -142 -153 -130 -119
rect -188 -187 -130 -153
rect -188 -221 -176 -187
rect -142 -221 -130 -187
rect -188 -255 -130 -221
rect -188 -289 -176 -255
rect -142 -289 -130 -255
rect -188 -323 -130 -289
rect -188 -357 -176 -323
rect -142 -357 -130 -323
rect -188 -391 -130 -357
rect -188 -425 -176 -391
rect -142 -425 -130 -391
rect -188 -459 -130 -425
rect -188 -493 -176 -459
rect -142 -493 -130 -459
rect -188 -527 -130 -493
rect -188 -561 -176 -527
rect -142 -561 -130 -527
rect -188 -595 -130 -561
rect -188 -629 -176 -595
rect -142 -629 -130 -595
rect -188 -663 -130 -629
rect -188 -697 -176 -663
rect -142 -697 -130 -663
rect -188 -731 -130 -697
rect -188 -765 -176 -731
rect -142 -765 -130 -731
rect -188 -799 -130 -765
rect -188 -833 -176 -799
rect -142 -833 -130 -799
rect -188 -867 -130 -833
rect -188 -901 -176 -867
rect -142 -901 -130 -867
rect -188 -935 -130 -901
rect -188 -969 -176 -935
rect -142 -969 -130 -935
rect -188 -1000 -130 -969
rect 130 969 188 1000
rect 130 935 142 969
rect 176 935 188 969
rect 130 901 188 935
rect 130 867 142 901
rect 176 867 188 901
rect 130 833 188 867
rect 130 799 142 833
rect 176 799 188 833
rect 130 765 188 799
rect 130 731 142 765
rect 176 731 188 765
rect 130 697 188 731
rect 130 663 142 697
rect 176 663 188 697
rect 130 629 188 663
rect 130 595 142 629
rect 176 595 188 629
rect 130 561 188 595
rect 130 527 142 561
rect 176 527 188 561
rect 130 493 188 527
rect 130 459 142 493
rect 176 459 188 493
rect 130 425 188 459
rect 130 391 142 425
rect 176 391 188 425
rect 130 357 188 391
rect 130 323 142 357
rect 176 323 188 357
rect 130 289 188 323
rect 130 255 142 289
rect 176 255 188 289
rect 130 221 188 255
rect 130 187 142 221
rect 176 187 188 221
rect 130 153 188 187
rect 130 119 142 153
rect 176 119 188 153
rect 130 85 188 119
rect 130 51 142 85
rect 176 51 188 85
rect 130 17 188 51
rect 130 -17 142 17
rect 176 -17 188 17
rect 130 -51 188 -17
rect 130 -85 142 -51
rect 176 -85 188 -51
rect 130 -119 188 -85
rect 130 -153 142 -119
rect 176 -153 188 -119
rect 130 -187 188 -153
rect 130 -221 142 -187
rect 176 -221 188 -187
rect 130 -255 188 -221
rect 130 -289 142 -255
rect 176 -289 188 -255
rect 130 -323 188 -289
rect 130 -357 142 -323
rect 176 -357 188 -323
rect 130 -391 188 -357
rect 130 -425 142 -391
rect 176 -425 188 -391
rect 130 -459 188 -425
rect 130 -493 142 -459
rect 176 -493 188 -459
rect 130 -527 188 -493
rect 130 -561 142 -527
rect 176 -561 188 -527
rect 130 -595 188 -561
rect 130 -629 142 -595
rect 176 -629 188 -595
rect 130 -663 188 -629
rect 130 -697 142 -663
rect 176 -697 188 -663
rect 130 -731 188 -697
rect 130 -765 142 -731
rect 176 -765 188 -731
rect 130 -799 188 -765
rect 130 -833 142 -799
rect 176 -833 188 -799
rect 130 -867 188 -833
rect 130 -901 142 -867
rect 176 -901 188 -867
rect 130 -935 188 -901
rect 130 -969 142 -935
rect 176 -969 188 -935
rect 130 -1000 188 -969
<< pdiffc >>
rect -176 935 -142 969
rect -176 867 -142 901
rect -176 799 -142 833
rect -176 731 -142 765
rect -176 663 -142 697
rect -176 595 -142 629
rect -176 527 -142 561
rect -176 459 -142 493
rect -176 391 -142 425
rect -176 323 -142 357
rect -176 255 -142 289
rect -176 187 -142 221
rect -176 119 -142 153
rect -176 51 -142 85
rect -176 -17 -142 17
rect -176 -85 -142 -51
rect -176 -153 -142 -119
rect -176 -221 -142 -187
rect -176 -289 -142 -255
rect -176 -357 -142 -323
rect -176 -425 -142 -391
rect -176 -493 -142 -459
rect -176 -561 -142 -527
rect -176 -629 -142 -595
rect -176 -697 -142 -663
rect -176 -765 -142 -731
rect -176 -833 -142 -799
rect -176 -901 -142 -867
rect -176 -969 -142 -935
rect 142 935 176 969
rect 142 867 176 901
rect 142 799 176 833
rect 142 731 176 765
rect 142 663 176 697
rect 142 595 176 629
rect 142 527 176 561
rect 142 459 176 493
rect 142 391 176 425
rect 142 323 176 357
rect 142 255 176 289
rect 142 187 176 221
rect 142 119 176 153
rect 142 51 176 85
rect 142 -17 176 17
rect 142 -85 176 -51
rect 142 -153 176 -119
rect 142 -221 176 -187
rect 142 -289 176 -255
rect 142 -357 176 -323
rect 142 -425 176 -391
rect 142 -493 176 -459
rect 142 -561 176 -527
rect 142 -629 176 -595
rect 142 -697 176 -663
rect 142 -765 176 -731
rect 142 -833 176 -799
rect 142 -901 176 -867
rect 142 -969 176 -935
<< nsubdiff >>
rect -290 1149 -187 1183
rect -153 1149 -119 1183
rect -85 1149 -51 1183
rect -17 1149 17 1183
rect 51 1149 85 1183
rect 119 1149 153 1183
rect 187 1149 290 1183
rect -290 1071 -256 1149
rect -290 1003 -256 1037
rect 256 1071 290 1149
rect 256 1003 290 1037
rect -290 935 -256 969
rect -290 867 -256 901
rect -290 799 -256 833
rect -290 731 -256 765
rect -290 663 -256 697
rect -290 595 -256 629
rect -290 527 -256 561
rect -290 459 -256 493
rect -290 391 -256 425
rect -290 323 -256 357
rect -290 255 -256 289
rect -290 187 -256 221
rect -290 119 -256 153
rect -290 51 -256 85
rect -290 -17 -256 17
rect -290 -85 -256 -51
rect -290 -153 -256 -119
rect -290 -221 -256 -187
rect -290 -289 -256 -255
rect -290 -357 -256 -323
rect -290 -425 -256 -391
rect -290 -493 -256 -459
rect -290 -561 -256 -527
rect -290 -629 -256 -595
rect -290 -697 -256 -663
rect -290 -765 -256 -731
rect -290 -833 -256 -799
rect -290 -901 -256 -867
rect -290 -969 -256 -935
rect 256 935 290 969
rect 256 867 290 901
rect 256 799 290 833
rect 256 731 290 765
rect 256 663 290 697
rect 256 595 290 629
rect 256 527 290 561
rect 256 459 290 493
rect 256 391 290 425
rect 256 323 290 357
rect 256 255 290 289
rect 256 187 290 221
rect 256 119 290 153
rect 256 51 290 85
rect 256 -17 290 17
rect 256 -85 290 -51
rect 256 -153 290 -119
rect 256 -221 290 -187
rect 256 -289 290 -255
rect 256 -357 290 -323
rect 256 -425 290 -391
rect 256 -493 290 -459
rect 256 -561 290 -527
rect 256 -629 290 -595
rect 256 -697 290 -663
rect 256 -765 290 -731
rect 256 -833 290 -799
rect 256 -901 290 -867
rect 256 -969 290 -935
rect -290 -1037 -256 -1003
rect -290 -1149 -256 -1071
rect 256 -1037 290 -1003
rect 256 -1149 290 -1071
rect -290 -1183 -187 -1149
rect -153 -1183 -119 -1149
rect -85 -1183 -51 -1149
rect -17 -1183 17 -1149
rect 51 -1183 85 -1149
rect 119 -1183 153 -1149
rect 187 -1183 290 -1149
<< nsubdiffcont >>
rect -187 1149 -153 1183
rect -119 1149 -85 1183
rect -51 1149 -17 1183
rect 17 1149 51 1183
rect 85 1149 119 1183
rect 153 1149 187 1183
rect -290 1037 -256 1071
rect -290 969 -256 1003
rect 256 1037 290 1071
rect -290 901 -256 935
rect -290 833 -256 867
rect -290 765 -256 799
rect -290 697 -256 731
rect -290 629 -256 663
rect -290 561 -256 595
rect -290 493 -256 527
rect -290 425 -256 459
rect -290 357 -256 391
rect -290 289 -256 323
rect -290 221 -256 255
rect -290 153 -256 187
rect -290 85 -256 119
rect -290 17 -256 51
rect -290 -51 -256 -17
rect -290 -119 -256 -85
rect -290 -187 -256 -153
rect -290 -255 -256 -221
rect -290 -323 -256 -289
rect -290 -391 -256 -357
rect -290 -459 -256 -425
rect -290 -527 -256 -493
rect -290 -595 -256 -561
rect -290 -663 -256 -629
rect -290 -731 -256 -697
rect -290 -799 -256 -765
rect -290 -867 -256 -833
rect -290 -935 -256 -901
rect -290 -1003 -256 -969
rect 256 969 290 1003
rect 256 901 290 935
rect 256 833 290 867
rect 256 765 290 799
rect 256 697 290 731
rect 256 629 290 663
rect 256 561 290 595
rect 256 493 290 527
rect 256 425 290 459
rect 256 357 290 391
rect 256 289 290 323
rect 256 221 290 255
rect 256 153 290 187
rect 256 85 290 119
rect 256 17 290 51
rect 256 -51 290 -17
rect 256 -119 290 -85
rect 256 -187 290 -153
rect 256 -255 290 -221
rect 256 -323 290 -289
rect 256 -391 290 -357
rect 256 -459 290 -425
rect 256 -527 290 -493
rect 256 -595 290 -561
rect 256 -663 290 -629
rect 256 -731 290 -697
rect 256 -799 290 -765
rect 256 -867 290 -833
rect 256 -935 290 -901
rect -290 -1071 -256 -1037
rect 256 -1003 290 -969
rect 256 -1071 290 -1037
rect -187 -1183 -153 -1149
rect -119 -1183 -85 -1149
rect -51 -1183 -17 -1149
rect 17 -1183 51 -1149
rect 85 -1183 119 -1149
rect 153 -1183 187 -1149
<< poly >>
rect -130 1081 130 1097
rect -130 1047 -85 1081
rect -51 1047 -17 1081
rect 17 1047 51 1081
rect 85 1047 130 1081
rect -130 1000 130 1047
rect -130 -1047 130 -1000
rect -130 -1081 -85 -1047
rect -51 -1081 -17 -1047
rect 17 -1081 51 -1047
rect 85 -1081 130 -1047
rect -130 -1097 130 -1081
<< polycont >>
rect -85 1047 -51 1081
rect -17 1047 17 1081
rect 51 1047 85 1081
rect -85 -1081 -51 -1047
rect -17 -1081 17 -1047
rect 51 -1081 85 -1047
<< locali >>
rect -290 1149 -187 1183
rect -153 1149 -119 1183
rect -85 1149 -51 1183
rect -17 1149 17 1183
rect 51 1149 85 1183
rect 119 1149 153 1183
rect 187 1149 290 1183
rect -290 1071 -256 1149
rect -130 1047 -89 1081
rect -51 1047 -17 1081
rect 17 1047 51 1081
rect 89 1047 130 1081
rect 256 1071 290 1149
rect -290 1003 -256 1037
rect -290 935 -256 969
rect -290 867 -256 901
rect -290 799 -256 833
rect -290 731 -256 765
rect -290 663 -256 697
rect -290 595 -256 629
rect -290 527 -256 561
rect -290 459 -256 493
rect -290 391 -256 425
rect -290 323 -256 357
rect -290 255 -256 289
rect -290 187 -256 221
rect -290 119 -256 153
rect -290 51 -256 85
rect -290 -17 -256 17
rect -290 -85 -256 -51
rect -290 -153 -256 -119
rect -290 -221 -256 -187
rect -290 -289 -256 -255
rect -290 -357 -256 -323
rect -290 -425 -256 -391
rect -290 -493 -256 -459
rect -290 -561 -256 -527
rect -290 -629 -256 -595
rect -290 -697 -256 -663
rect -290 -765 -256 -731
rect -290 -833 -256 -799
rect -290 -901 -256 -867
rect -290 -969 -256 -935
rect -290 -1037 -256 -1003
rect -176 969 -142 1004
rect -176 901 -142 919
rect -176 833 -142 847
rect -176 765 -142 775
rect -176 697 -142 703
rect -176 629 -142 631
rect -176 593 -142 595
rect -176 521 -142 527
rect -176 449 -142 459
rect -176 377 -142 391
rect -176 305 -142 323
rect -176 233 -142 255
rect -176 161 -142 187
rect -176 89 -142 119
rect -176 17 -142 51
rect -176 -51 -142 -17
rect -176 -119 -142 -89
rect -176 -187 -142 -161
rect -176 -255 -142 -233
rect -176 -323 -142 -305
rect -176 -391 -142 -377
rect -176 -459 -142 -449
rect -176 -527 -142 -521
rect -176 -595 -142 -593
rect -176 -631 -142 -629
rect -176 -703 -142 -697
rect -176 -775 -142 -765
rect -176 -847 -142 -833
rect -176 -919 -142 -901
rect -176 -1004 -142 -969
rect 142 969 176 1004
rect 142 901 176 919
rect 142 833 176 847
rect 142 765 176 775
rect 142 697 176 703
rect 142 629 176 631
rect 142 593 176 595
rect 142 521 176 527
rect 142 449 176 459
rect 142 377 176 391
rect 142 305 176 323
rect 142 233 176 255
rect 142 161 176 187
rect 142 89 176 119
rect 142 17 176 51
rect 142 -51 176 -17
rect 142 -119 176 -89
rect 142 -187 176 -161
rect 142 -255 176 -233
rect 142 -323 176 -305
rect 142 -391 176 -377
rect 142 -459 176 -449
rect 142 -527 176 -521
rect 142 -595 176 -593
rect 142 -631 176 -629
rect 142 -703 176 -697
rect 142 -775 176 -765
rect 142 -847 176 -833
rect 142 -919 176 -901
rect 142 -1004 176 -969
rect 256 1003 290 1037
rect 256 935 290 969
rect 256 867 290 901
rect 256 799 290 833
rect 256 731 290 765
rect 256 663 290 697
rect 256 595 290 629
rect 256 527 290 561
rect 256 459 290 493
rect 256 391 290 425
rect 256 323 290 357
rect 256 255 290 289
rect 256 187 290 221
rect 256 119 290 153
rect 256 51 290 85
rect 256 -17 290 17
rect 256 -85 290 -51
rect 256 -153 290 -119
rect 256 -221 290 -187
rect 256 -289 290 -255
rect 256 -357 290 -323
rect 256 -425 290 -391
rect 256 -493 290 -459
rect 256 -561 290 -527
rect 256 -629 290 -595
rect 256 -697 290 -663
rect 256 -765 290 -731
rect 256 -833 290 -799
rect 256 -901 290 -867
rect 256 -969 290 -935
rect 256 -1037 290 -1003
rect -290 -1149 -256 -1071
rect -130 -1081 -89 -1047
rect -51 -1081 -17 -1047
rect 17 -1081 51 -1047
rect 89 -1081 130 -1047
rect 256 -1149 290 -1071
rect -290 -1183 -187 -1149
rect -153 -1183 -119 -1149
rect -85 -1183 -51 -1149
rect -17 -1183 17 -1149
rect 51 -1183 85 -1149
rect 119 -1183 153 -1149
rect 187 -1183 290 -1149
<< viali >>
rect -89 1047 -85 1081
rect -85 1047 -55 1081
rect -17 1047 17 1081
rect 55 1047 85 1081
rect 85 1047 89 1081
rect -176 935 -142 953
rect -176 919 -142 935
rect -176 867 -142 881
rect -176 847 -142 867
rect -176 799 -142 809
rect -176 775 -142 799
rect -176 731 -142 737
rect -176 703 -142 731
rect -176 663 -142 665
rect -176 631 -142 663
rect -176 561 -142 593
rect -176 559 -142 561
rect -176 493 -142 521
rect -176 487 -142 493
rect -176 425 -142 449
rect -176 415 -142 425
rect -176 357 -142 377
rect -176 343 -142 357
rect -176 289 -142 305
rect -176 271 -142 289
rect -176 221 -142 233
rect -176 199 -142 221
rect -176 153 -142 161
rect -176 127 -142 153
rect -176 85 -142 89
rect -176 55 -142 85
rect -176 -17 -142 17
rect -176 -85 -142 -55
rect -176 -89 -142 -85
rect -176 -153 -142 -127
rect -176 -161 -142 -153
rect -176 -221 -142 -199
rect -176 -233 -142 -221
rect -176 -289 -142 -271
rect -176 -305 -142 -289
rect -176 -357 -142 -343
rect -176 -377 -142 -357
rect -176 -425 -142 -415
rect -176 -449 -142 -425
rect -176 -493 -142 -487
rect -176 -521 -142 -493
rect -176 -561 -142 -559
rect -176 -593 -142 -561
rect -176 -663 -142 -631
rect -176 -665 -142 -663
rect -176 -731 -142 -703
rect -176 -737 -142 -731
rect -176 -799 -142 -775
rect -176 -809 -142 -799
rect -176 -867 -142 -847
rect -176 -881 -142 -867
rect -176 -935 -142 -919
rect -176 -953 -142 -935
rect 142 935 176 953
rect 142 919 176 935
rect 142 867 176 881
rect 142 847 176 867
rect 142 799 176 809
rect 142 775 176 799
rect 142 731 176 737
rect 142 703 176 731
rect 142 663 176 665
rect 142 631 176 663
rect 142 561 176 593
rect 142 559 176 561
rect 142 493 176 521
rect 142 487 176 493
rect 142 425 176 449
rect 142 415 176 425
rect 142 357 176 377
rect 142 343 176 357
rect 142 289 176 305
rect 142 271 176 289
rect 142 221 176 233
rect 142 199 176 221
rect 142 153 176 161
rect 142 127 176 153
rect 142 85 176 89
rect 142 55 176 85
rect 142 -17 176 17
rect 142 -85 176 -55
rect 142 -89 176 -85
rect 142 -153 176 -127
rect 142 -161 176 -153
rect 142 -221 176 -199
rect 142 -233 176 -221
rect 142 -289 176 -271
rect 142 -305 176 -289
rect 142 -357 176 -343
rect 142 -377 176 -357
rect 142 -425 176 -415
rect 142 -449 176 -425
rect 142 -493 176 -487
rect 142 -521 176 -493
rect 142 -561 176 -559
rect 142 -593 176 -561
rect 142 -663 176 -631
rect 142 -665 176 -663
rect 142 -731 176 -703
rect 142 -737 176 -731
rect 142 -799 176 -775
rect 142 -809 176 -799
rect 142 -867 176 -847
rect 142 -881 176 -867
rect 142 -935 176 -919
rect 142 -953 176 -935
rect -89 -1081 -85 -1047
rect -85 -1081 -55 -1047
rect -17 -1081 17 -1047
rect 55 -1081 85 -1047
rect 85 -1081 89 -1047
<< metal1 >>
rect -126 1081 126 1087
rect -126 1047 -89 1081
rect -55 1047 -17 1081
rect 17 1047 55 1081
rect 89 1047 126 1081
rect -126 1041 126 1047
rect -182 953 -136 1000
rect -182 919 -176 953
rect -142 919 -136 953
rect -182 881 -136 919
rect -182 847 -176 881
rect -142 847 -136 881
rect -182 809 -136 847
rect -182 775 -176 809
rect -142 775 -136 809
rect -182 737 -136 775
rect -182 703 -176 737
rect -142 703 -136 737
rect -182 665 -136 703
rect -182 631 -176 665
rect -142 631 -136 665
rect -182 593 -136 631
rect -182 559 -176 593
rect -142 559 -136 593
rect -182 521 -136 559
rect -182 487 -176 521
rect -142 487 -136 521
rect -182 449 -136 487
rect -182 415 -176 449
rect -142 415 -136 449
rect -182 377 -136 415
rect -182 343 -176 377
rect -142 343 -136 377
rect -182 305 -136 343
rect -182 271 -176 305
rect -142 271 -136 305
rect -182 233 -136 271
rect -182 199 -176 233
rect -142 199 -136 233
rect -182 161 -136 199
rect -182 127 -176 161
rect -142 127 -136 161
rect -182 89 -136 127
rect -182 55 -176 89
rect -142 55 -136 89
rect -182 17 -136 55
rect -182 -17 -176 17
rect -142 -17 -136 17
rect -182 -55 -136 -17
rect -182 -89 -176 -55
rect -142 -89 -136 -55
rect -182 -127 -136 -89
rect -182 -161 -176 -127
rect -142 -161 -136 -127
rect -182 -199 -136 -161
rect -182 -233 -176 -199
rect -142 -233 -136 -199
rect -182 -271 -136 -233
rect -182 -305 -176 -271
rect -142 -305 -136 -271
rect -182 -343 -136 -305
rect -182 -377 -176 -343
rect -142 -377 -136 -343
rect -182 -415 -136 -377
rect -182 -449 -176 -415
rect -142 -449 -136 -415
rect -182 -487 -136 -449
rect -182 -521 -176 -487
rect -142 -521 -136 -487
rect -182 -559 -136 -521
rect -182 -593 -176 -559
rect -142 -593 -136 -559
rect -182 -631 -136 -593
rect -182 -665 -176 -631
rect -142 -665 -136 -631
rect -182 -703 -136 -665
rect -182 -737 -176 -703
rect -142 -737 -136 -703
rect -182 -775 -136 -737
rect -182 -809 -176 -775
rect -142 -809 -136 -775
rect -182 -847 -136 -809
rect -182 -881 -176 -847
rect -142 -881 -136 -847
rect -182 -919 -136 -881
rect -182 -953 -176 -919
rect -142 -953 -136 -919
rect -182 -1000 -136 -953
rect 136 953 182 1000
rect 136 919 142 953
rect 176 919 182 953
rect 136 881 182 919
rect 136 847 142 881
rect 176 847 182 881
rect 136 809 182 847
rect 136 775 142 809
rect 176 775 182 809
rect 136 737 182 775
rect 136 703 142 737
rect 176 703 182 737
rect 136 665 182 703
rect 136 631 142 665
rect 176 631 182 665
rect 136 593 182 631
rect 136 559 142 593
rect 176 559 182 593
rect 136 521 182 559
rect 136 487 142 521
rect 176 487 182 521
rect 136 449 182 487
rect 136 415 142 449
rect 176 415 182 449
rect 136 377 182 415
rect 136 343 142 377
rect 176 343 182 377
rect 136 305 182 343
rect 136 271 142 305
rect 176 271 182 305
rect 136 233 182 271
rect 136 199 142 233
rect 176 199 182 233
rect 136 161 182 199
rect 136 127 142 161
rect 176 127 182 161
rect 136 89 182 127
rect 136 55 142 89
rect 176 55 182 89
rect 136 17 182 55
rect 136 -17 142 17
rect 176 -17 182 17
rect 136 -55 182 -17
rect 136 -89 142 -55
rect 176 -89 182 -55
rect 136 -127 182 -89
rect 136 -161 142 -127
rect 176 -161 182 -127
rect 136 -199 182 -161
rect 136 -233 142 -199
rect 176 -233 182 -199
rect 136 -271 182 -233
rect 136 -305 142 -271
rect 176 -305 182 -271
rect 136 -343 182 -305
rect 136 -377 142 -343
rect 176 -377 182 -343
rect 136 -415 182 -377
rect 136 -449 142 -415
rect 176 -449 182 -415
rect 136 -487 182 -449
rect 136 -521 142 -487
rect 176 -521 182 -487
rect 136 -559 182 -521
rect 136 -593 142 -559
rect 176 -593 182 -559
rect 136 -631 182 -593
rect 136 -665 142 -631
rect 176 -665 182 -631
rect 136 -703 182 -665
rect 136 -737 142 -703
rect 176 -737 182 -703
rect 136 -775 182 -737
rect 136 -809 142 -775
rect 176 -809 182 -775
rect 136 -847 182 -809
rect 136 -881 142 -847
rect 176 -881 182 -847
rect 136 -919 182 -881
rect 136 -953 142 -919
rect 176 -953 182 -919
rect 136 -1000 182 -953
rect -126 -1047 126 -1041
rect -126 -1081 -89 -1047
rect -55 -1081 -17 -1047
rect 17 -1081 55 -1047
rect 89 -1081 126 -1047
rect -126 -1087 126 -1081
<< properties >>
string FIXED_BBOX -273 -1166 273 1166
<< end >>
