magic
tech sky130A
magscale 1 2
timestamp 1716990733
<< pwell >>
rect -686 -257 686 257
<< nmos >>
rect -500 -57 500 57
<< ndiff >>
rect -558 17 -500 57
rect -558 -17 -546 17
rect -512 -17 -500 17
rect -558 -57 -500 -17
rect 500 17 558 57
rect 500 -17 512 17
rect 546 -17 558 17
rect 500 -57 558 -17
<< ndiffc >>
rect -546 -17 -512 17
rect 512 -17 546 17
<< psubdiff >>
rect -660 197 -561 231
rect -527 197 -493 231
rect -459 197 -425 231
rect -391 197 -357 231
rect -323 197 -289 231
rect -255 197 -221 231
rect -187 197 -153 231
rect -119 197 -85 231
rect -51 197 -17 231
rect 17 197 51 231
rect 85 197 119 231
rect 153 197 187 231
rect 221 197 255 231
rect 289 197 323 231
rect 357 197 391 231
rect 425 197 459 231
rect 493 197 527 231
rect 561 197 660 231
rect -660 119 -626 197
rect -660 51 -626 85
rect 626 119 660 197
rect -660 -17 -626 17
rect -660 -85 -626 -51
rect 626 51 660 85
rect 626 -17 660 17
rect -660 -197 -626 -119
rect 626 -85 660 -51
rect 626 -197 660 -119
rect -660 -231 -561 -197
rect -527 -231 -493 -197
rect -459 -231 -425 -197
rect -391 -231 -357 -197
rect -323 -231 -289 -197
rect -255 -231 -221 -197
rect -187 -231 -153 -197
rect -119 -231 -85 -197
rect -51 -231 -17 -197
rect 17 -231 51 -197
rect 85 -231 119 -197
rect 153 -231 187 -197
rect 221 -231 255 -197
rect 289 -231 323 -197
rect 357 -231 391 -197
rect 425 -231 459 -197
rect 493 -231 527 -197
rect 561 -231 660 -197
<< psubdiffcont >>
rect -561 197 -527 231
rect -493 197 -459 231
rect -425 197 -391 231
rect -357 197 -323 231
rect -289 197 -255 231
rect -221 197 -187 231
rect -153 197 -119 231
rect -85 197 -51 231
rect -17 197 17 231
rect 51 197 85 231
rect 119 197 153 231
rect 187 197 221 231
rect 255 197 289 231
rect 323 197 357 231
rect 391 197 425 231
rect 459 197 493 231
rect 527 197 561 231
rect -660 85 -626 119
rect 626 85 660 119
rect -660 17 -626 51
rect -660 -51 -626 -17
rect 626 17 660 51
rect 626 -51 660 -17
rect -660 -119 -626 -85
rect 626 -119 660 -85
rect -561 -231 -527 -197
rect -493 -231 -459 -197
rect -425 -231 -391 -197
rect -357 -231 -323 -197
rect -289 -231 -255 -197
rect -221 -231 -187 -197
rect -153 -231 -119 -197
rect -85 -231 -51 -197
rect -17 -231 17 -197
rect 51 -231 85 -197
rect 119 -231 153 -197
rect 187 -231 221 -197
rect 255 -231 289 -197
rect 323 -231 357 -197
rect 391 -231 425 -197
rect 459 -231 493 -197
rect 527 -231 561 -197
<< poly >>
rect -500 129 500 145
rect -500 95 -459 129
rect -425 95 -391 129
rect -357 95 -323 129
rect -289 95 -255 129
rect -221 95 -187 129
rect -153 95 -119 129
rect -85 95 -51 129
rect -17 95 17 129
rect 51 95 85 129
rect 119 95 153 129
rect 187 95 221 129
rect 255 95 289 129
rect 323 95 357 129
rect 391 95 425 129
rect 459 95 500 129
rect -500 57 500 95
rect -500 -95 500 -57
rect -500 -129 -459 -95
rect -425 -129 -391 -95
rect -357 -129 -323 -95
rect -289 -129 -255 -95
rect -221 -129 -187 -95
rect -153 -129 -119 -95
rect -85 -129 -51 -95
rect -17 -129 17 -95
rect 51 -129 85 -95
rect 119 -129 153 -95
rect 187 -129 221 -95
rect 255 -129 289 -95
rect 323 -129 357 -95
rect 391 -129 425 -95
rect 459 -129 500 -95
rect -500 -145 500 -129
<< polycont >>
rect -459 95 -425 129
rect -391 95 -357 129
rect -323 95 -289 129
rect -255 95 -221 129
rect -187 95 -153 129
rect -119 95 -85 129
rect -51 95 -17 129
rect 17 95 51 129
rect 85 95 119 129
rect 153 95 187 129
rect 221 95 255 129
rect 289 95 323 129
rect 357 95 391 129
rect 425 95 459 129
rect -459 -129 -425 -95
rect -391 -129 -357 -95
rect -323 -129 -289 -95
rect -255 -129 -221 -95
rect -187 -129 -153 -95
rect -119 -129 -85 -95
rect -51 -129 -17 -95
rect 17 -129 51 -95
rect 85 -129 119 -95
rect 153 -129 187 -95
rect 221 -129 255 -95
rect 289 -129 323 -95
rect 357 -129 391 -95
rect 425 -129 459 -95
<< locali >>
rect -660 197 -561 231
rect -527 197 -493 231
rect -459 197 -425 231
rect -391 197 -357 231
rect -323 197 -289 231
rect -255 197 -221 231
rect -187 197 -153 231
rect -119 197 -85 231
rect -51 197 -17 231
rect 17 197 51 231
rect 85 197 119 231
rect 153 197 187 231
rect 221 197 255 231
rect 289 197 323 231
rect 357 197 391 231
rect 425 197 459 231
rect 493 197 527 231
rect 561 197 660 231
rect -660 119 -626 197
rect -500 95 -459 129
rect -415 95 -391 129
rect -343 95 -323 129
rect -271 95 -255 129
rect -199 95 -187 129
rect -127 95 -119 129
rect -55 95 -51 129
rect 51 95 55 129
rect 119 95 127 129
rect 187 95 199 129
rect 255 95 271 129
rect 323 95 343 129
rect 391 95 415 129
rect 459 95 500 129
rect 626 119 660 197
rect -660 51 -626 85
rect -660 -17 -626 17
rect -660 -85 -626 -51
rect -546 17 -512 61
rect -546 -61 -512 -17
rect 512 17 546 61
rect 512 -61 546 -17
rect 626 51 660 85
rect 626 -17 660 17
rect 626 -85 660 -51
rect -660 -197 -626 -119
rect -500 -129 -459 -95
rect -415 -129 -391 -95
rect -343 -129 -323 -95
rect -271 -129 -255 -95
rect -199 -129 -187 -95
rect -127 -129 -119 -95
rect -55 -129 -51 -95
rect 51 -129 55 -95
rect 119 -129 127 -95
rect 187 -129 199 -95
rect 255 -129 271 -95
rect 323 -129 343 -95
rect 391 -129 415 -95
rect 459 -129 500 -95
rect 626 -197 660 -119
rect -660 -231 -561 -197
rect -527 -231 -493 -197
rect -459 -231 -425 -197
rect -391 -231 -357 -197
rect -323 -231 -289 -197
rect -255 -231 -221 -197
rect -187 -231 -153 -197
rect -119 -231 -85 -197
rect -51 -231 -17 -197
rect 17 -231 51 -197
rect 85 -231 119 -197
rect 153 -231 187 -197
rect 221 -231 255 -197
rect 289 -231 323 -197
rect 357 -231 391 -197
rect 425 -231 459 -197
rect 493 -231 527 -197
rect 561 -231 660 -197
<< viali >>
rect -449 95 -425 129
rect -425 95 -415 129
rect -377 95 -357 129
rect -357 95 -343 129
rect -305 95 -289 129
rect -289 95 -271 129
rect -233 95 -221 129
rect -221 95 -199 129
rect -161 95 -153 129
rect -153 95 -127 129
rect -89 95 -85 129
rect -85 95 -55 129
rect -17 95 17 129
rect 55 95 85 129
rect 85 95 89 129
rect 127 95 153 129
rect 153 95 161 129
rect 199 95 221 129
rect 221 95 233 129
rect 271 95 289 129
rect 289 95 305 129
rect 343 95 357 129
rect 357 95 377 129
rect 415 95 425 129
rect 425 95 449 129
rect -546 -17 -512 17
rect 512 -17 546 17
rect -449 -129 -425 -95
rect -425 -129 -415 -95
rect -377 -129 -357 -95
rect -357 -129 -343 -95
rect -305 -129 -289 -95
rect -289 -129 -271 -95
rect -233 -129 -221 -95
rect -221 -129 -199 -95
rect -161 -129 -153 -95
rect -153 -129 -127 -95
rect -89 -129 -85 -95
rect -85 -129 -55 -95
rect -17 -129 17 -95
rect 55 -129 85 -95
rect 85 -129 89 -95
rect 127 -129 153 -95
rect 153 -129 161 -95
rect 199 -129 221 -95
rect 221 -129 233 -95
rect 271 -129 289 -95
rect 289 -129 305 -95
rect 343 -129 357 -95
rect 357 -129 377 -95
rect 415 -129 425 -95
rect 425 -129 449 -95
<< metal1 >>
rect -496 129 496 135
rect -496 95 -449 129
rect -415 95 -377 129
rect -343 95 -305 129
rect -271 95 -233 129
rect -199 95 -161 129
rect -127 95 -89 129
rect -55 95 -17 129
rect 17 95 55 129
rect 89 95 127 129
rect 161 95 199 129
rect 233 95 271 129
rect 305 95 343 129
rect 377 95 415 129
rect 449 95 496 129
rect -496 89 496 95
rect -552 17 -506 57
rect -552 -17 -546 17
rect -512 -17 -506 17
rect -552 -57 -506 -17
rect 506 17 552 57
rect 506 -17 512 17
rect 546 -17 552 17
rect 506 -57 552 -17
rect -496 -95 496 -89
rect -496 -129 -449 -95
rect -415 -129 -377 -95
rect -343 -129 -305 -95
rect -271 -129 -233 -95
rect -199 -129 -161 -95
rect -127 -129 -89 -95
rect -55 -129 -17 -95
rect 17 -129 55 -95
rect 89 -129 127 -95
rect 161 -129 199 -95
rect 233 -129 271 -95
rect 305 -129 343 -95
rect 377 -129 415 -95
rect 449 -129 496 -95
rect -496 -135 496 -129
<< properties >>
string FIXED_BBOX -643 -214 643 214
<< end >>
