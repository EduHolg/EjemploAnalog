MACRO sky130_fd_pr__pfet_01v8_NXK9QA
  CLASS BLOCK ;
  FOREIGN sky130_fd_pr__pfet_01v8_NXK9QA ;
  ORIGIN 2.215 2.330 ;
  SIZE 4.430 BY 4.660 ;
  OBS
      LAYER nwell ;
        RECT -2.480 -2.595 2.480 2.595 ;
      LAYER li1 ;
        RECT -2.300 2.245 2.300 2.415 ;
        RECT -2.300 -2.245 -2.130 2.245 ;
        RECT -1.500 1.735 1.500 1.905 ;
        RECT -1.730 -1.520 -1.560 1.520 ;
        RECT 1.560 -1.520 1.730 1.520 ;
        RECT -1.500 -1.905 1.500 -1.735 ;
        RECT 2.130 -2.245 2.300 2.245 ;
        RECT -2.300 -2.415 2.300 -2.245 ;
      LAYER mcon ;
        RECT -1.345 1.735 -1.175 1.905 ;
        RECT -0.985 1.735 -0.815 1.905 ;
        RECT -0.625 1.735 -0.455 1.905 ;
        RECT -0.265 1.735 -0.095 1.905 ;
        RECT 0.095 1.735 0.265 1.905 ;
        RECT 0.455 1.735 0.625 1.905 ;
        RECT 0.815 1.735 0.985 1.905 ;
        RECT 1.175 1.735 1.345 1.905 ;
        RECT -1.730 1.175 -1.560 1.345 ;
        RECT -1.730 0.815 -1.560 0.985 ;
        RECT -1.730 0.455 -1.560 0.625 ;
        RECT -1.730 0.095 -1.560 0.265 ;
        RECT -1.730 -0.265 -1.560 -0.095 ;
        RECT -1.730 -0.625 -1.560 -0.455 ;
        RECT -1.730 -0.985 -1.560 -0.815 ;
        RECT -1.730 -1.345 -1.560 -1.175 ;
        RECT 1.560 1.175 1.730 1.345 ;
        RECT 1.560 0.815 1.730 0.985 ;
        RECT 1.560 0.455 1.730 0.625 ;
        RECT 1.560 0.095 1.730 0.265 ;
        RECT 1.560 -0.265 1.730 -0.095 ;
        RECT 1.560 -0.625 1.730 -0.455 ;
        RECT 1.560 -0.985 1.730 -0.815 ;
        RECT 1.560 -1.345 1.730 -1.175 ;
        RECT -1.345 -1.905 -1.175 -1.735 ;
        RECT -0.985 -1.905 -0.815 -1.735 ;
        RECT -0.625 -1.905 -0.455 -1.735 ;
        RECT -0.265 -1.905 -0.095 -1.735 ;
        RECT 0.095 -1.905 0.265 -1.735 ;
        RECT 0.455 -1.905 0.625 -1.735 ;
        RECT 0.815 -1.905 0.985 -1.735 ;
        RECT 1.175 -1.905 1.345 -1.735 ;
      LAYER met1 ;
        RECT -1.480 1.705 1.480 1.935 ;
        RECT -1.760 -1.500 -1.530 1.500 ;
        RECT 1.530 -1.500 1.760 1.500 ;
        RECT -1.480 -1.935 1.480 -1.705 ;
  END
END sky130_fd_pr__pfet_01v8_NXK9QA
END LIBRARY

